library ieee;
-- muss noch fertig schreiben!
